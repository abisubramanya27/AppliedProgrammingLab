.circuit
R1 N002 N003 1e3
V1 N001 GND ac 5 0
C1 N002 N001 1
L1 N003 GND 1e-6
.end
.ac 1e3