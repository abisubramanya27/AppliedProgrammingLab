.circuit
V1 N001 GND ac 1 0
R1 N002 N001 4.5e3
R2 GND N004 4e3
L1 N002 N003 80.96e-6
L2 N003 N004 80.96e-6
C1 N003 GND 2.485e-12
.end
.ac 1e3